/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HD__UDP_PWRGOOD_L_PP_PG_S_TB_V
`define SKY130_FD_SC_HD__UDP_PWRGOOD_L_PP_PG_S_TB_V

/**

 *   UDP_OUT :=x when VPWR!=1 or VGND!=0
 *   UDP_OUT :=UDP_IN when VPWR==1 and VGND==0
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none


module top();

    // Inputs are registered
    reg UDP_IN;
    reg VPWR;
    reg VGND;
    reg SLEEP;

    // Outputs are wires
    wire UDP_OUT;

    initial
    begin
        // Initial state is x for all inputs.
        SLEEP  = 1'bX;
        UDP_IN = 1'bX;
        VGND   = 1'bX;
        VPWR   = 1'bX;

        #20   SLEEP  = 1'b0;
        #40   UDP_IN = 1'b0;
        #60   VGND   = 1'b0;
        #80   VPWR   = 1'b0;
        #100  SLEEP  = 1'b1;
        #120  UDP_IN = 1'b1;
        #140  VGND   = 1'b1;
        #160  VPWR   = 1'b1;
        #180  SLEEP  = 1'b0;
        #200  UDP_IN = 1'b0;
        #220  VGND   = 1'b0;
        #240  VPWR   = 1'b0;
        #260  VPWR   = 1'b1;
        #280  VGND   = 1'b1;
        #300  UDP_IN = 1'b1;
        #320  SLEEP  = 1'b1;
        #340  VPWR   = 1'bx;
        #360  VGND   = 1'bx;
        #380  UDP_IN = 1'bx;
        #400  SLEEP  = 1'bx;
    end

    sky130_fd_sc_hd__udp_pwrgood$l_pp$PG$S dut (.UDP_IN(UDP_IN), .VPWR(VPWR), .VGND(VGND), .SLEEP(SLEEP), .UDP_OUT(UDP_OUT));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HD__UDP_PWRGOOD_L_PP_PG_S_TB_V
